
module alu_sim (
    input  logic clk_i,
    input  logic rst_ni,
    input  logic rxd_i,
    output logic txd_o
);

alu alu (.*);

endmodule
