package dv_pkg;

import config_pkg::*;

// put DV params/tasks/functions here

endpackage